package gcd_pkg;
    `include "gcd_packet.sv"
	`include "generator.sv"
    `include "calc_gcd.sv"
    `include "driver.sv"
	`include "scoreboard.sv"
    `include "monitor.sv"
endpackage